`include "defines.v"

module mainControl (
    input 
);
    
endmodule